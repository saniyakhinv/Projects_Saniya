library ieee;
use ieee.std_logic_1164.all;
package Flipflops is
	component dff_set is port(D,clock,set:in std_logic;Q:out std_logic);
	end component dff_set;
	component dff_reset is port(D,clock,reset:in std_logic:='0';Q:out std_logic:='0');
	end component dff_reset;
end package Flipflops;

--D flip flop with set

library ieee;
use ieee.std_logic_1164.all;
entity dff_set is port(D,clock,set:in std_logic; Q:out std_logic);
end entity dff_set;
architecture behav of dff_set is
begin
	dff_set_proc: process (clock,set)
	begin
		if(set='1')then -- set implies flip flip output logic high
		Q <='1' ; -- write the flip flop output when set
		elsif (clock'event and (clock='1')) then
		Q <=D ; -- write flip flop output when not set
		end if ;
	end process dff_set_proc;
end behav;

--D flip flop with reset
library ieee;
use ieee.std_logic_1164.all;
entity dff_reset is port(D,clock,reset:in std_logic:='0'; Q:out std_logic:='0');
end entity dff_reset;
architecture behav of dff_reset is
begin
	dff_reset_proc: process (clock,reset)
	begin
		if(reset='1')then -- reset implies flip flip output logic low
		Q <='0'; -- write the flip flop output when reset
		elsif (falling_edge(clock)) then
		Q <=D ; -- write flip flop output when not reset
		
		end if ;
	end process dff_reset_proc;
end behav;